`timescale 1ns / 1ps
module InstructionMemory(PC_Address, Instruction);
input [31:0] PC_Address;
output [31:0] Instruction;
/*
parameter InstMem_size = 512;
reg [31:0] instruction [InstMem_size-1:0];
*/
assign Instruction =	
    (PC_Address[9:2] == 8'd0)?32'h2004003c:
    (PC_Address[9:2] == 8'd1)?32'h20050000:
    (PC_Address[9:2] == 8'd2)?32'h20060004:
    (PC_Address[9:2] == 8'd3)?32'h20070190:
    (PC_Address[9:2] == 8'd4)?32'h20080000:
    (PC_Address[9:2] == 8'd5)?32'h20100000:
    (PC_Address[9:2] == 8'd6)?32'h00865022:
    (PC_Address[9:2] == 8'd7)?32'h214a0001:
    (PC_Address[9:2] == 8'd8)?32'h20cb0001:
    (PC_Address[9:2] == 8'd9)?32'h110a000f:
    (PC_Address[9:2] == 8'd10)?32'h20090000:
    (PC_Address[9:2] == 8'd11)?32'h112b0008:
    (PC_Address[9:2] == 8'd12)?32'h01096020:
    (PC_Address[9:2] == 8'd13)?32'h01856820:
    (PC_Address[9:2] == 8'd14)?32'h81ae0000:
    (PC_Address[9:2] == 8'd15)?32'h01276020:
    (PC_Address[9:2] == 8'd16)?32'h818d0000:
    (PC_Address[9:2] == 8'd17)?32'h21290001:
    (PC_Address[9:2] == 8'd18)?32'h15ae0001:
    (PC_Address[9:2] == 8'd19)?32'h0810000b:
    (PC_Address[9:2] == 8'd20)?32'h21080001:
    (PC_Address[9:2] == 8'd21)?32'h112b0001:
    (PC_Address[9:2] == 8'd22)?32'h08100009:
    (PC_Address[9:2] == 8'd23)?32'h22100001:
    (PC_Address[9:2] == 8'd24)?32'h08100009:
    (PC_Address[9:2] == 8'd25)?32'h00101020:
    (PC_Address[9:2] == 8'd26)?32'h20100000:
    (PC_Address[9:2] == 8'd27)?32'h00104302:
    (PC_Address[9:2] == 8'd28)?32'h31080003:
    (PC_Address[9:2] == 8'd29)?32'h20090000:
    (PC_Address[9:2] == 8'd30)?32'h11090006:
    (PC_Address[9:2] == 8'd31)?32'h21290001:
    (PC_Address[9:2] == 8'd32)?32'h11090007:
    (PC_Address[9:2] == 8'd33)?32'h21290001:
    (PC_Address[9:2] == 8'd34)?32'h11090009:
    (PC_Address[9:2] == 8'd35)?32'h21290001:
    (PC_Address[9:2] == 8'd36)?32'h1109000b:
    (PC_Address[9:2] == 8'd37)?32'h20110100:
    (PC_Address[9:2] == 8'd38)?32'h304a000f:
    (PC_Address[9:2] == 8'd39)?32'h08100033:
    (PC_Address[9:2] == 8'd40)?32'h20110200:
    (PC_Address[9:2] == 8'd41)?32'h304a00f0:
    (PC_Address[9:2] == 8'd42)?32'h000a5102:
    (PC_Address[9:2] == 8'd43)?32'h08100033:
    (PC_Address[9:2] == 8'd44)?32'h20110400:
    (PC_Address[9:2] == 8'd45)?32'h304a0f00:
    (PC_Address[9:2] == 8'd46)?32'h000a5202:
    (PC_Address[9:2] == 8'd47)?32'h08100033:
    (PC_Address[9:2] == 8'd48)?32'h20110800:
    (PC_Address[9:2] == 8'd49)?32'h304af000:
    (PC_Address[9:2] == 8'd50)?32'h000a5302:
    (PC_Address[9:2] == 8'd51)?32'h20090000:
    (PC_Address[9:2] == 8'd52)?32'h1149001e:
    (PC_Address[9:2] == 8'd53)?32'h21290001:
    (PC_Address[9:2] == 8'd54)?32'h1149001e:
    (PC_Address[9:2] == 8'd55)?32'h21290001:
    (PC_Address[9:2] == 8'd56)?32'h1149001e:
    (PC_Address[9:2] == 8'd57)?32'h21290001:
    (PC_Address[9:2] == 8'd58)?32'h1149001e:
    (PC_Address[9:2] == 8'd59)?32'h21290001:
    (PC_Address[9:2] == 8'd60)?32'h1149001e:
    (PC_Address[9:2] == 8'd61)?32'h21290001:
    (PC_Address[9:2] == 8'd62)?32'h1149001e:
    (PC_Address[9:2] == 8'd63)?32'h21290001:
    (PC_Address[9:2] == 8'd64)?32'h1149001e:
    (PC_Address[9:2] == 8'd65)?32'h21290001:
    (PC_Address[9:2] == 8'd66)?32'h1149001e:
    (PC_Address[9:2] == 8'd67)?32'h21290001:
    (PC_Address[9:2] == 8'd68)?32'h1149001e:
    (PC_Address[9:2] == 8'd69)?32'h21290001:
    (PC_Address[9:2] == 8'd70)?32'h1149001e:
    (PC_Address[9:2] == 8'd71)?32'h21290001:
    (PC_Address[9:2] == 8'd72)?32'h1149001e:
    (PC_Address[9:2] == 8'd73)?32'h21290001:
    (PC_Address[9:2] == 8'd74)?32'h1149001e:
    (PC_Address[9:2] == 8'd75)?32'h21290001:
    (PC_Address[9:2] == 8'd76)?32'h1149001e:
    (PC_Address[9:2] == 8'd77)?32'h21290001:
    (PC_Address[9:2] == 8'd78)?32'h1149001e:
    (PC_Address[9:2] == 8'd79)?32'h21290001:
    (PC_Address[9:2] == 8'd80)?32'h1149001e:
    (PC_Address[9:2] == 8'd81)?32'h21290001:
    (PC_Address[9:2] == 8'd82)?32'h1149001e:
    (PC_Address[9:2] == 8'd83)?32'h200b003f:
    (PC_Address[9:2] == 8'd84)?32'h08100072:
    (PC_Address[9:2] == 8'd85)?32'h200b0006:
    (PC_Address[9:2] == 8'd86)?32'h08100072:
    (PC_Address[9:2] == 8'd87)?32'h200b005b:
    (PC_Address[9:2] == 8'd88)?32'h08100072:
    (PC_Address[9:2] == 8'd89)?32'h200b004f:
    (PC_Address[9:2] == 8'd90)?32'h08100072:
    (PC_Address[9:2] == 8'd91)?32'h200b0066:
    (PC_Address[9:2] == 8'd92)?32'h08100072:
    (PC_Address[9:2] == 8'd93)?32'h200b006d:
    (PC_Address[9:2] == 8'd94)?32'h08100072:
    (PC_Address[9:2] == 8'd95)?32'h200b007d:
    (PC_Address[9:2] == 8'd96)?32'h08100072:
    (PC_Address[9:2] == 8'd97)?32'h200b0007:
    (PC_Address[9:2] == 8'd98)?32'h08100072:
    (PC_Address[9:2] == 8'd99)?32'h200b007f:
    (PC_Address[9:2] == 8'd100)?32'h08100072:
    (PC_Address[9:2] == 8'd101)?32'h200b006f:
    (PC_Address[9:2] == 8'd102)?32'h08100072:
    (PC_Address[9:2] == 8'd103)?32'h200b0077:
    (PC_Address[9:2] == 8'd104)?32'h08100072:
    (PC_Address[9:2] == 8'd105)?32'h200b007c:
    (PC_Address[9:2] == 8'd106)?32'h08100072:
    (PC_Address[9:2] == 8'd107)?32'h200b0039:
    (PC_Address[9:2] == 8'd108)?32'h08100072:
    (PC_Address[9:2] == 8'd109)?32'h200b005e:
    (PC_Address[9:2] == 8'd110)?32'h08100072:
    (PC_Address[9:2] == 8'd111)?32'h200b0079:
    (PC_Address[9:2] == 8'd112)?32'h08100072:
    (PC_Address[9:2] == 8'd113)?32'h200b0071:
    (PC_Address[9:2] == 8'd114)?32'h022b9020:
    (PC_Address[9:2] == 8'd115)?32'h200c4000:
    (PC_Address[9:2] == 8'd116)?32'h000c6400:
    (PC_Address[9:2] == 8'd117)?32'h218c0010:
    (PC_Address[9:2] == 8'd118)?32'had920000:
    (PC_Address[9:2] == 8'd119)?32'h22100001:
    (PC_Address[9:2] == 8'd120)?32'h0810001b:
  32'h00000000;

endmodule
